library verilog;
use verilog.vl_types.all;
entity BUF_X16 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end BUF_X16;
