library verilog;
use verilog.vl_types.all;
entity seq43 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end seq43;
