library verilog;
use verilog.vl_types.all;
entity ANTENNA_X1 is
    port(
        A               : in     vl_logic
    );
end ANTENNA_X1;
