library verilog;
use verilog.vl_types.all;
entity FILLCELL_X8 is
end FILLCELL_X8;
