library verilog;
use verilog.vl_types.all;
entity CLKBUF_X2 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end CLKBUF_X2;
