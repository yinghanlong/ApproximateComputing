library verilog;
use verilog.vl_types.all;
entity FILLCELL_X4 is
end FILLCELL_X4;
