library verilog;
use verilog.vl_types.all;
entity OAI211_X4 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end OAI211_X4;
