library verilog;
use verilog.vl_types.all;
entity FILLCELL_X2 is
end FILLCELL_X2;
