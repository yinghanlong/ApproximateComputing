library verilog;
use verilog.vl_types.all;
entity FILLCELL_X1 is
end FILLCELL_X1;
