library verilog;
use verilog.vl_types.all;
entity FILLCELL_X16 is
end FILLCELL_X16;
