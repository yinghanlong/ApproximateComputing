library verilog;
use verilog.vl_types.all;
entity test_fixture is
end test_fixture;
