library verilog;
use verilog.vl_types.all;
entity AOI22_X4 is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end AOI22_X4;
