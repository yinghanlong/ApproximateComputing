library verilog;
use verilog.vl_types.all;
entity FILLCELL_X32 is
end FILLCELL_X32;
